module enc2freq (
    input logic cw, ccw,        // outputs from lab 2 encoder module
    output logic [31:10] freq,  // desired frequency
    input logic reset_n, clk);  // reset and clock

    

endmodule