module tonegen
    #( parameter FCLK )
    ( input logic [31:0] freq,